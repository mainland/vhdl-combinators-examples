library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.lava.all;
use work.all;
entity incrementer is
  port(clk : in std_logic;
       in_x : in std_logic_vector(15 downto 0);
       reset : in std_logic;
       in_valid : in std_logic;
       out_ready : in std_logic;
       out_valid : out std_logic;
       in_ready : out std_logic;
       out_x : out std_logic_vector(15 downto 0));
end entity incrementer;
architecture str of incrementer is
  signal sig_237_o0 : std_logic_vector(15 downto 0);
  signal sig_238_o0 : std_logic_vector(15 downto 0);
  signal sig_235_o0 : std_logic;
  signal sig_236_o0 : std_logic;
  signal sig_2_o0 : std_logic;
  signal sig_3_o0 : std_logic;
  signal sig_4_o0 : std_logic_vector(17 downto 0);
  signal sig_234_o0 : std_logic;
  signal sig_233_o0 : std_logic;
  signal sig_5_o0 : std_logic_vector(15 downto 0);
  signal sig_6_o0 : std_logic_vector(16 downto 0);
  signal sig_232_o0 : std_logic_vector(15 downto 0);
  signal sig_7_o0 : std_logic;
  signal sig_8_o0 : std_logic_vector(16 downto 0);
  signal sig_143_o0 : std_logic_vector(15 downto 0);
  type sig_144_o0_type is array (31 downto 0) of std_logic_vector(15 downto 0);
  signal sig_144_o0 : sig_144_o0_type;
  type sig_145_o0_type is array (31 downto 0) of std_logic_vector(15 downto 0);
  signal sig_145_o0 : sig_145_o0_type;
  type sig_146_o0_type is array (31 downto 0) of std_logic_vector(15 downto 0);
  signal sig_146_o0 : sig_146_o0_type;
  signal sig_227_o0 : std_logic_vector(15 downto 0);
  signal sig_230_o0 : std_logic_vector(15 downto 0);
  signal sig_231_o0 : std_logic_vector(15 downto 0);
  signal sig_228_o0 : std_logic_vector(15 downto 0);
  signal sig_229_o0 : std_logic_vector(15 downto 0);
  signal sig_222_o0 : std_logic_vector(15 downto 0);
  signal sig_225_o0 : std_logic_vector(15 downto 0);
  signal sig_226_o0 : std_logic_vector(15 downto 0);
  signal sig_223_o0 : std_logic_vector(15 downto 0);
  signal sig_224_o0 : std_logic_vector(15 downto 0);
  signal sig_217_o0 : std_logic_vector(15 downto 0);
  signal sig_220_o0 : std_logic_vector(15 downto 0);
  signal sig_221_o0 : std_logic_vector(15 downto 0);
  signal sig_218_o0 : std_logic_vector(15 downto 0);
  signal sig_219_o0 : std_logic_vector(15 downto 0);
  signal sig_212_o0 : std_logic_vector(15 downto 0);
  signal sig_215_o0 : std_logic_vector(15 downto 0);
  signal sig_216_o0 : std_logic_vector(15 downto 0);
  signal sig_213_o0 : std_logic_vector(15 downto 0);
  signal sig_214_o0 : std_logic_vector(15 downto 0);
  signal sig_207_o0 : std_logic_vector(15 downto 0);
  signal sig_210_o0 : std_logic_vector(15 downto 0);
  signal sig_211_o0 : std_logic_vector(15 downto 0);
  signal sig_208_o0 : std_logic_vector(15 downto 0);
  signal sig_209_o0 : std_logic_vector(15 downto 0);
  signal sig_202_o0 : std_logic_vector(15 downto 0);
  signal sig_205_o0 : std_logic_vector(15 downto 0);
  signal sig_206_o0 : std_logic_vector(15 downto 0);
  signal sig_203_o0 : std_logic_vector(15 downto 0);
  signal sig_204_o0 : std_logic_vector(15 downto 0);
  signal sig_197_o0 : std_logic_vector(15 downto 0);
  signal sig_200_o0 : std_logic_vector(15 downto 0);
  signal sig_201_o0 : std_logic_vector(15 downto 0);
  signal sig_198_o0 : std_logic_vector(15 downto 0);
  signal sig_199_o0 : std_logic_vector(15 downto 0);
  signal sig_192_o0 : std_logic_vector(15 downto 0);
  signal sig_195_o0 : std_logic_vector(15 downto 0);
  signal sig_196_o0 : std_logic_vector(15 downto 0);
  signal sig_193_o0 : std_logic_vector(15 downto 0);
  signal sig_194_o0 : std_logic_vector(15 downto 0);
  signal sig_187_o0 : std_logic_vector(15 downto 0);
  signal sig_190_o0 : std_logic_vector(15 downto 0);
  signal sig_191_o0 : std_logic_vector(15 downto 0);
  signal sig_188_o0 : std_logic_vector(15 downto 0);
  signal sig_189_o0 : std_logic_vector(15 downto 0);
  signal sig_182_o0 : std_logic_vector(15 downto 0);
  signal sig_185_o0 : std_logic_vector(15 downto 0);
  signal sig_186_o0 : std_logic_vector(15 downto 0);
  signal sig_183_o0 : std_logic_vector(15 downto 0);
  signal sig_184_o0 : std_logic_vector(15 downto 0);
  signal sig_177_o0 : std_logic_vector(15 downto 0);
  signal sig_180_o0 : std_logic_vector(15 downto 0);
  signal sig_181_o0 : std_logic_vector(15 downto 0);
  signal sig_178_o0 : std_logic_vector(15 downto 0);
  signal sig_179_o0 : std_logic_vector(15 downto 0);
  signal sig_172_o0 : std_logic_vector(15 downto 0);
  signal sig_175_o0 : std_logic_vector(15 downto 0);
  signal sig_176_o0 : std_logic_vector(15 downto 0);
  signal sig_173_o0 : std_logic_vector(15 downto 0);
  signal sig_174_o0 : std_logic_vector(15 downto 0);
  signal sig_167_o0 : std_logic_vector(15 downto 0);
  signal sig_170_o0 : std_logic_vector(15 downto 0);
  signal sig_171_o0 : std_logic_vector(15 downto 0);
  signal sig_168_o0 : std_logic_vector(15 downto 0);
  signal sig_169_o0 : std_logic_vector(15 downto 0);
  signal sig_162_o0 : std_logic_vector(15 downto 0);
  signal sig_165_o0 : std_logic_vector(15 downto 0);
  signal sig_166_o0 : std_logic_vector(15 downto 0);
  signal sig_163_o0 : std_logic_vector(15 downto 0);
  signal sig_164_o0 : std_logic_vector(15 downto 0);
  signal sig_157_o0 : std_logic_vector(15 downto 0);
  signal sig_160_o0 : std_logic_vector(15 downto 0);
  signal sig_161_o0 : std_logic_vector(15 downto 0);
  signal sig_158_o0 : std_logic_vector(15 downto 0);
  signal sig_159_o0 : std_logic_vector(15 downto 0);
  signal sig_152_o0 : std_logic_vector(15 downto 0);
  signal sig_155_o0 : std_logic_vector(15 downto 0);
  signal sig_156_o0 : std_logic_vector(15 downto 0);
  signal sig_153_o0 : std_logic_vector(15 downto 0);
  signal sig_154_o0 : std_logic_vector(15 downto 0);
  signal sig_147_o0 : std_logic_vector(15 downto 0);
  signal sig_150_o0 : std_logic_vector(15 downto 0);
  signal sig_151_o0 : std_logic_vector(15 downto 0);
  signal sig_148_o0 : std_logic_vector(15 downto 0);
  signal sig_149_o0 : std_logic_vector(15 downto 0);
  signal sig_9_o0 : std_logic;
  type sig_10_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_10_o0 : sig_10_o0_type;
  type sig_11_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_11_o0 : sig_11_o0_type;
  type sig_142_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_142_o0 : sig_142_o0_type;
  type sig_13_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_13_o0 : sig_13_o0_type;
  type sig_16_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_16_o0 : sig_16_o0_type;
  signal sig_138_o0 : std_logic;
  signal sig_140_o0 : std_logic;
  signal sig_141_o0 : std_logic;
  signal sig_139_o0 : std_logic;
  signal sig_135_o0 : std_logic;
  signal sig_136_o0 : std_logic;
  signal sig_137_o0 : std_logic;
  signal sig_132_o0 : std_logic;
  signal sig_133_o0 : std_logic;
  signal sig_134_o0 : std_logic;
  signal sig_129_o0 : std_logic;
  signal sig_130_o0 : std_logic;
  signal sig_131_o0 : std_logic;
  signal sig_126_o0 : std_logic;
  signal sig_127_o0 : std_logic;
  signal sig_128_o0 : std_logic;
  signal sig_123_o0 : std_logic;
  signal sig_124_o0 : std_logic;
  signal sig_125_o0 : std_logic;
  signal sig_120_o0 : std_logic;
  signal sig_121_o0 : std_logic;
  signal sig_122_o0 : std_logic;
  signal sig_117_o0 : std_logic;
  signal sig_118_o0 : std_logic;
  signal sig_119_o0 : std_logic;
  signal sig_114_o0 : std_logic;
  signal sig_115_o0 : std_logic;
  signal sig_116_o0 : std_logic;
  signal sig_111_o0 : std_logic;
  signal sig_112_o0 : std_logic;
  signal sig_113_o0 : std_logic;
  signal sig_108_o0 : std_logic;
  signal sig_109_o0 : std_logic;
  signal sig_110_o0 : std_logic;
  signal sig_105_o0 : std_logic;
  signal sig_106_o0 : std_logic;
  signal sig_107_o0 : std_logic;
  signal sig_102_o0 : std_logic;
  signal sig_103_o0 : std_logic;
  signal sig_104_o0 : std_logic;
  signal sig_99_o0 : std_logic;
  signal sig_100_o0 : std_logic;
  signal sig_101_o0 : std_logic;
  signal sig_96_o0 : std_logic;
  signal sig_97_o0 : std_logic;
  signal sig_98_o0 : std_logic;
  signal sig_93_o0 : std_logic;
  signal sig_94_o0 : std_logic;
  signal sig_95_o0 : std_logic;
  signal sig_17_o0 : std_logic;
  signal sig_92_o0 : std_logic;
  signal sig_90_o0 : std_logic;
  signal sig_91_o0 : std_logic;
  signal sig_18_o0 : std_logic;
  type sig_19_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_19_o0 : sig_19_o0_type;
  type sig_89_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_89_o0 : sig_89_o0_type;
  type sig_20_o0_type is array (31 downto 0) of std_logic_vector(0 downto 0);
  signal sig_20_o0 : sig_20_o0_type;
  signal sig_81_o0 : std_logic;
  signal sig_87_o0 : std_logic;
  signal sig_88_o0 : std_logic;
  signal sig_82_o0 : std_logic;
  signal sig_83_o0 : std_logic_vector(17 downto 0);
  signal sig_86_o0 : std_logic;
  signal sig_85_o0 : std_logic;
  signal sig_84_o0 : std_logic_vector(15 downto 0);
  signal sig_77_o0 : std_logic;
  signal sig_79_o0 : std_logic;
  signal sig_80_o0 : std_logic;
  signal sig_78_o0 : std_logic;
  signal sig_73_o0 : std_logic;
  signal sig_75_o0 : std_logic;
  signal sig_76_o0 : std_logic;
  signal sig_74_o0 : std_logic;
  signal sig_69_o0 : std_logic;
  signal sig_71_o0 : std_logic;
  signal sig_72_o0 : std_logic;
  signal sig_70_o0 : std_logic;
  signal sig_65_o0 : std_logic;
  signal sig_67_o0 : std_logic;
  signal sig_68_o0 : std_logic;
  signal sig_66_o0 : std_logic;
  signal sig_61_o0 : std_logic;
  signal sig_63_o0 : std_logic;
  signal sig_64_o0 : std_logic;
  signal sig_62_o0 : std_logic;
  signal sig_57_o0 : std_logic;
  signal sig_59_o0 : std_logic;
  signal sig_60_o0 : std_logic;
  signal sig_58_o0 : std_logic;
  signal sig_53_o0 : std_logic;
  signal sig_55_o0 : std_logic;
  signal sig_56_o0 : std_logic;
  signal sig_54_o0 : std_logic;
  signal sig_49_o0 : std_logic;
  signal sig_51_o0 : std_logic;
  signal sig_52_o0 : std_logic;
  signal sig_50_o0 : std_logic;
  signal sig_45_o0 : std_logic;
  signal sig_47_o0 : std_logic;
  signal sig_48_o0 : std_logic;
  signal sig_46_o0 : std_logic;
  signal sig_41_o0 : std_logic;
  signal sig_43_o0 : std_logic;
  signal sig_44_o0 : std_logic;
  signal sig_42_o0 : std_logic;
  signal sig_37_o0 : std_logic;
  signal sig_39_o0 : std_logic;
  signal sig_40_o0 : std_logic;
  signal sig_38_o0 : std_logic;
  signal sig_33_o0 : std_logic;
  signal sig_35_o0 : std_logic;
  signal sig_36_o0 : std_logic;
  signal sig_34_o0 : std_logic;
  signal sig_29_o0 : std_logic;
  signal sig_31_o0 : std_logic;
  signal sig_32_o0 : std_logic;
  signal sig_30_o0 : std_logic;
  signal sig_25_o0 : std_logic;
  signal sig_27_o0 : std_logic;
  signal sig_28_o0 : std_logic;
  signal sig_26_o0 : std_logic;
  signal sig_21_o0 : std_logic;
  signal sig_23_o0 : std_logic;
  signal sig_24_o0 : std_logic;
  signal sig_22_o0 : std_logic;
  signal sig_14_o0 : std_logic;
  signal sig_15_o0 : std_logic;
  signal sig_12_o0 : std_logic;
begin
  sig_237_o0 <= sig_238_o0;
  sig_238_o0 <= sig_4_o0(15 downto 0);
  sig_235_o0 <= sig_236_o0;
  sig_236_o0 <= sig_4_o0(17);
  sig_2_o0 <= sig_3_o0;
  sig_3_o0 <= sig_4_o0(16);
  -- [("i0",16U,(5).o0),("i1",B,(233).o0),("i2",B,(234).o0)];
  sig_4_o0 <= sig_234_o0 & sig_233_o0 & sig_5_o0;
  sig_234_o0 <= lava_to_std_logic(sig_19_o0(0));
  sig_233_o0 <= sig_6_o0(0);
  sig_5_o0 <= sig_6_o0(16 downto 1);
  -- [("i0",B,(7).o0),("i1",16U,(232).o0)];
  sig_6_o0 <= sig_232_o0 & sig_7_o0;
  sig_232_o0 <= sig_8_o0(16 downto 1);
  sig_7_o0 <= sig_8_o0(0);
  -- [("i0",B,(9).o0),("i1",16U,(143).o0)];
  sig_8_o0 <= sig_143_o0 & sig_9_o0;
  sig_143_o0 <= sig_144_o0(15);
  proc255 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_144_o0(0) <= sig_145_o0(0);
        sig_144_o0(1) <= sig_145_o0(1);
        sig_144_o0(2) <= sig_145_o0(2);
        sig_144_o0(3) <= sig_145_o0(3);
        sig_144_o0(4) <= sig_145_o0(4);
        sig_144_o0(5) <= sig_145_o0(5);
        sig_144_o0(6) <= sig_145_o0(6);
        sig_144_o0(7) <= sig_145_o0(7);
        sig_144_o0(8) <= sig_145_o0(8);
        sig_144_o0(9) <= sig_145_o0(9);
        sig_144_o0(10) <= sig_145_o0(10);
        sig_144_o0(11) <= sig_145_o0(11);
        sig_144_o0(12) <= sig_145_o0(12);
        sig_144_o0(13) <= sig_145_o0(13);
        sig_144_o0(14) <= sig_145_o0(14);
        sig_144_o0(15) <= sig_145_o0(15);
        sig_144_o0(16) <= sig_145_o0(16);
      end if;
    end if;
  end process proc255;
  sig_145_o0(0) <= sig_146_o0(0) when (sig_14_o0 = '1') else
                   sig_144_o0(0);
  sig_145_o0(1) <= sig_146_o0(1) when (sig_14_o0 = '1') else
                   sig_144_o0(1);
  sig_145_o0(2) <= sig_146_o0(2) when (sig_14_o0 = '1') else
                   sig_144_o0(2);
  sig_145_o0(3) <= sig_146_o0(3) when (sig_14_o0 = '1') else
                   sig_144_o0(3);
  sig_145_o0(4) <= sig_146_o0(4) when (sig_14_o0 = '1') else
                   sig_144_o0(4);
  sig_145_o0(5) <= sig_146_o0(5) when (sig_14_o0 = '1') else
                   sig_144_o0(5);
  sig_145_o0(6) <= sig_146_o0(6) when (sig_14_o0 = '1') else
                   sig_144_o0(6);
  sig_145_o0(7) <= sig_146_o0(7) when (sig_14_o0 = '1') else
                   sig_144_o0(7);
  sig_145_o0(8) <= sig_146_o0(8) when (sig_14_o0 = '1') else
                   sig_144_o0(8);
  sig_145_o0(9) <= sig_146_o0(9) when (sig_14_o0 = '1') else
                   sig_144_o0(9);
  sig_145_o0(10) <= sig_146_o0(10) when (sig_14_o0 = '1') else
                    sig_144_o0(10);
  sig_145_o0(11) <= sig_146_o0(11) when (sig_14_o0 = '1') else
                    sig_144_o0(11);
  sig_145_o0(12) <= sig_146_o0(12) when (sig_14_o0 = '1') else
                    sig_144_o0(12);
  sig_145_o0(13) <= sig_146_o0(13) when (sig_14_o0 = '1') else
                    sig_144_o0(13);
  sig_145_o0(14) <= sig_146_o0(14) when (sig_14_o0 = '1') else
                    sig_144_o0(14);
  sig_145_o0(15) <= sig_146_o0(15) when (sig_14_o0 = '1') else
                    sig_144_o0(15);
  sig_145_o0(16) <= sig_146_o0(16) when (sig_14_o0 = '1') else
                    sig_144_o0(16);
  sig_146_o0(0) <= sig_147_o0;
  sig_146_o0(1) <= sig_152_o0;
  sig_146_o0(2) <= sig_157_o0;
  sig_146_o0(3) <= sig_162_o0;
  sig_146_o0(4) <= sig_167_o0;
  sig_146_o0(5) <= sig_172_o0;
  sig_146_o0(6) <= sig_177_o0;
  sig_146_o0(7) <= sig_182_o0;
  sig_146_o0(8) <= sig_187_o0;
  sig_146_o0(9) <= sig_192_o0;
  sig_146_o0(10) <= sig_197_o0;
  sig_146_o0(11) <= sig_202_o0;
  sig_146_o0(12) <= sig_207_o0;
  sig_146_o0(13) <= sig_212_o0;
  sig_146_o0(14) <= sig_217_o0;
  sig_146_o0(15) <= sig_222_o0;
  sig_146_o0(16) <= sig_227_o0;
  sig_227_o0 <= sig_230_o0 when (sig_139_o0 = '1') else
                sig_228_o0;
  sig_230_o0 <= std_logic_vector((unsigned(sig_231_o0) + to_unsigned(1,
                                                                     16)));
  sig_231_o0 <= sig_144_o0(15);
  proc293 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_228_o0 <= sig_229_o0;
      end if;
    end if;
  end process proc293;
  sig_229_o0 <= sig_145_o0(16);
  sig_222_o0 <= sig_225_o0 when (sig_78_o0 = '1') else
                sig_223_o0;
  sig_225_o0 <= std_logic_vector((unsigned(sig_226_o0) + to_unsigned(1,
                                                                     16)));
  sig_226_o0 <= sig_144_o0(14);
  proc298 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_223_o0 <= sig_224_o0;
      end if;
    end if;
  end process proc298;
  sig_224_o0 <= sig_145_o0(15);
  sig_217_o0 <= sig_220_o0 when (sig_74_o0 = '1') else
                sig_218_o0;
  sig_220_o0 <= std_logic_vector((unsigned(sig_221_o0) + to_unsigned(1,
                                                                     16)));
  sig_221_o0 <= sig_144_o0(13);
  proc303 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_218_o0 <= sig_219_o0;
      end if;
    end if;
  end process proc303;
  sig_219_o0 <= sig_145_o0(14);
  sig_212_o0 <= sig_215_o0 when (sig_70_o0 = '1') else
                sig_213_o0;
  sig_215_o0 <= std_logic_vector((unsigned(sig_216_o0) + to_unsigned(1,
                                                                     16)));
  sig_216_o0 <= sig_144_o0(12);
  proc308 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_213_o0 <= sig_214_o0;
      end if;
    end if;
  end process proc308;
  sig_214_o0 <= sig_145_o0(13);
  sig_207_o0 <= sig_210_o0 when (sig_66_o0 = '1') else
                sig_208_o0;
  sig_210_o0 <= std_logic_vector((unsigned(sig_211_o0) + to_unsigned(1,
                                                                     16)));
  sig_211_o0 <= sig_144_o0(11);
  proc313 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_208_o0 <= sig_209_o0;
      end if;
    end if;
  end process proc313;
  sig_209_o0 <= sig_145_o0(12);
  sig_202_o0 <= sig_205_o0 when (sig_62_o0 = '1') else
                sig_203_o0;
  sig_205_o0 <= std_logic_vector((unsigned(sig_206_o0) + to_unsigned(1,
                                                                     16)));
  sig_206_o0 <= sig_144_o0(10);
  proc318 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_203_o0 <= sig_204_o0;
      end if;
    end if;
  end process proc318;
  sig_204_o0 <= sig_145_o0(11);
  sig_197_o0 <= sig_200_o0 when (sig_58_o0 = '1') else
                sig_198_o0;
  sig_200_o0 <= std_logic_vector((unsigned(sig_201_o0) + to_unsigned(1,
                                                                     16)));
  sig_201_o0 <= sig_144_o0(9);
  proc323 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_198_o0 <= sig_199_o0;
      end if;
    end if;
  end process proc323;
  sig_199_o0 <= sig_145_o0(10);
  sig_192_o0 <= sig_195_o0 when (sig_54_o0 = '1') else
                sig_193_o0;
  sig_195_o0 <= std_logic_vector((unsigned(sig_196_o0) + to_unsigned(1,
                                                                     16)));
  sig_196_o0 <= sig_144_o0(8);
  proc328 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_193_o0 <= sig_194_o0;
      end if;
    end if;
  end process proc328;
  sig_194_o0 <= sig_145_o0(9);
  sig_187_o0 <= sig_190_o0 when (sig_50_o0 = '1') else
                sig_188_o0;
  sig_190_o0 <= std_logic_vector((unsigned(sig_191_o0) + to_unsigned(1,
                                                                     16)));
  sig_191_o0 <= sig_144_o0(7);
  proc333 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_188_o0 <= sig_189_o0;
      end if;
    end if;
  end process proc333;
  sig_189_o0 <= sig_145_o0(8);
  sig_182_o0 <= sig_185_o0 when (sig_46_o0 = '1') else
                sig_183_o0;
  sig_185_o0 <= std_logic_vector((unsigned(sig_186_o0) + to_unsigned(1,
                                                                     16)));
  sig_186_o0 <= sig_144_o0(6);
  proc338 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_183_o0 <= sig_184_o0;
      end if;
    end if;
  end process proc338;
  sig_184_o0 <= sig_145_o0(7);
  sig_177_o0 <= sig_180_o0 when (sig_42_o0 = '1') else
                sig_178_o0;
  sig_180_o0 <= std_logic_vector((unsigned(sig_181_o0) + to_unsigned(1,
                                                                     16)));
  sig_181_o0 <= sig_144_o0(5);
  proc343 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_178_o0 <= sig_179_o0;
      end if;
    end if;
  end process proc343;
  sig_179_o0 <= sig_145_o0(6);
  sig_172_o0 <= sig_175_o0 when (sig_38_o0 = '1') else
                sig_173_o0;
  sig_175_o0 <= std_logic_vector((unsigned(sig_176_o0) + to_unsigned(1,
                                                                     16)));
  sig_176_o0 <= sig_144_o0(4);
  proc348 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_173_o0 <= sig_174_o0;
      end if;
    end if;
  end process proc348;
  sig_174_o0 <= sig_145_o0(5);
  sig_167_o0 <= sig_170_o0 when (sig_34_o0 = '1') else
                sig_168_o0;
  sig_170_o0 <= std_logic_vector((unsigned(sig_171_o0) + to_unsigned(1,
                                                                     16)));
  sig_171_o0 <= sig_144_o0(3);
  proc353 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_168_o0 <= sig_169_o0;
      end if;
    end if;
  end process proc353;
  sig_169_o0 <= sig_145_o0(4);
  sig_162_o0 <= sig_165_o0 when (sig_30_o0 = '1') else
                sig_163_o0;
  sig_165_o0 <= std_logic_vector((unsigned(sig_166_o0) + to_unsigned(1,
                                                                     16)));
  sig_166_o0 <= sig_144_o0(2);
  proc358 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_163_o0 <= sig_164_o0;
      end if;
    end if;
  end process proc358;
  sig_164_o0 <= sig_145_o0(3);
  sig_157_o0 <= sig_160_o0 when (sig_26_o0 = '1') else
                sig_158_o0;
  sig_160_o0 <= std_logic_vector((unsigned(sig_161_o0) + to_unsigned(1,
                                                                     16)));
  sig_161_o0 <= sig_144_o0(1);
  proc363 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_158_o0 <= sig_159_o0;
      end if;
    end if;
  end process proc363;
  sig_159_o0 <= sig_145_o0(2);
  sig_152_o0 <= sig_155_o0 when (sig_22_o0 = '1') else
                sig_153_o0;
  sig_155_o0 <= std_logic_vector((unsigned(sig_156_o0) + to_unsigned(1,
                                                                     16)));
  sig_156_o0 <= sig_144_o0(0);
  proc368 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_153_o0 <= sig_154_o0;
      end if;
    end if;
  end process proc368;
  sig_154_o0 <= sig_145_o0(1);
  sig_147_o0 <= sig_150_o0 when (sig_18_o0 = '1') else
                sig_148_o0;
  sig_150_o0 <= std_logic_vector((unsigned(sig_151_o0) + to_unsigned(1,
                                                                     16)));
  sig_151_o0 <= sig_83_o0(15 downto 0);
  proc373 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_148_o0 <= sig_149_o0;
      end if;
    end if;
  end process proc373;
  sig_149_o0 <= sig_145_o0(0);
  sig_9_o0 <= lava_to_std_logic(sig_10_o0(15));
  proc376 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_10_o0(0) <= sig_11_o0(0);
        sig_10_o0(1) <= sig_11_o0(1);
        sig_10_o0(2) <= sig_11_o0(2);
        sig_10_o0(3) <= sig_11_o0(3);
        sig_10_o0(4) <= sig_11_o0(4);
        sig_10_o0(5) <= sig_11_o0(5);
        sig_10_o0(6) <= sig_11_o0(6);
        sig_10_o0(7) <= sig_11_o0(7);
        sig_10_o0(8) <= sig_11_o0(8);
        sig_10_o0(9) <= sig_11_o0(9);
        sig_10_o0(10) <= sig_11_o0(10);
        sig_10_o0(11) <= sig_11_o0(11);
        sig_10_o0(12) <= sig_11_o0(12);
        sig_10_o0(13) <= sig_11_o0(13);
        sig_10_o0(14) <= sig_11_o0(14);
        sig_10_o0(15) <= sig_11_o0(15);
        sig_10_o0(16) <= sig_11_o0(16);
      end if;
    end if;
  end process proc376;
  sig_11_o0(0) <= sig_142_o0(0) when (sig_12_o0 = '1') else
                  sig_13_o0(0);
  sig_11_o0(1) <= sig_142_o0(1) when (sig_12_o0 = '1') else
                  sig_13_o0(1);
  sig_11_o0(2) <= sig_142_o0(2) when (sig_12_o0 = '1') else
                  sig_13_o0(2);
  sig_11_o0(3) <= sig_142_o0(3) when (sig_12_o0 = '1') else
                  sig_13_o0(3);
  sig_11_o0(4) <= sig_142_o0(4) when (sig_12_o0 = '1') else
                  sig_13_o0(4);
  sig_11_o0(5) <= sig_142_o0(5) when (sig_12_o0 = '1') else
                  sig_13_o0(5);
  sig_11_o0(6) <= sig_142_o0(6) when (sig_12_o0 = '1') else
                  sig_13_o0(6);
  sig_11_o0(7) <= sig_142_o0(7) when (sig_12_o0 = '1') else
                  sig_13_o0(7);
  sig_11_o0(8) <= sig_142_o0(8) when (sig_12_o0 = '1') else
                  sig_13_o0(8);
  sig_11_o0(9) <= sig_142_o0(9) when (sig_12_o0 = '1') else
                  sig_13_o0(9);
  sig_11_o0(10) <= sig_142_o0(10) when (sig_12_o0 = '1') else
                   sig_13_o0(10);
  sig_11_o0(11) <= sig_142_o0(11) when (sig_12_o0 = '1') else
                   sig_13_o0(11);
  sig_11_o0(12) <= sig_142_o0(12) when (sig_12_o0 = '1') else
                   sig_13_o0(12);
  sig_11_o0(13) <= sig_142_o0(13) when (sig_12_o0 = '1') else
                   sig_13_o0(13);
  sig_11_o0(14) <= sig_142_o0(14) when (sig_12_o0 = '1') else
                   sig_13_o0(14);
  sig_11_o0(15) <= sig_142_o0(15) when (sig_12_o0 = '1') else
                   sig_13_o0(15);
  sig_11_o0(16) <= sig_142_o0(16) when (sig_12_o0 = '1') else
                   sig_13_o0(16);
  sig_142_o0(0) <= "" & '0';
  sig_142_o0(1) <= "" & '0';
  sig_142_o0(2) <= "" & '0';
  sig_142_o0(3) <= "" & '0';
  sig_142_o0(4) <= "" & '0';
  sig_142_o0(5) <= "" & '0';
  sig_142_o0(6) <= "" & '0';
  sig_142_o0(7) <= "" & '0';
  sig_142_o0(8) <= "" & '0';
  sig_142_o0(9) <= "" & '0';
  sig_142_o0(10) <= "" & '0';
  sig_142_o0(11) <= "" & '0';
  sig_142_o0(12) <= "" & '0';
  sig_142_o0(13) <= "" & '0';
  sig_142_o0(14) <= "" & '0';
  sig_142_o0(15) <= "" & '0';
  sig_142_o0(16) <= "" & '0';
  sig_13_o0(0) <= sig_16_o0(0) when (sig_14_o0 = '1') else
                  sig_10_o0(0);
  sig_13_o0(1) <= sig_16_o0(1) when (sig_14_o0 = '1') else
                  sig_10_o0(1);
  sig_13_o0(2) <= sig_16_o0(2) when (sig_14_o0 = '1') else
                  sig_10_o0(2);
  sig_13_o0(3) <= sig_16_o0(3) when (sig_14_o0 = '1') else
                  sig_10_o0(3);
  sig_13_o0(4) <= sig_16_o0(4) when (sig_14_o0 = '1') else
                  sig_10_o0(4);
  sig_13_o0(5) <= sig_16_o0(5) when (sig_14_o0 = '1') else
                  sig_10_o0(5);
  sig_13_o0(6) <= sig_16_o0(6) when (sig_14_o0 = '1') else
                  sig_10_o0(6);
  sig_13_o0(7) <= sig_16_o0(7) when (sig_14_o0 = '1') else
                  sig_10_o0(7);
  sig_13_o0(8) <= sig_16_o0(8) when (sig_14_o0 = '1') else
                  sig_10_o0(8);
  sig_13_o0(9) <= sig_16_o0(9) when (sig_14_o0 = '1') else
                  sig_10_o0(9);
  sig_13_o0(10) <= sig_16_o0(10) when (sig_14_o0 = '1') else
                   sig_10_o0(10);
  sig_13_o0(11) <= sig_16_o0(11) when (sig_14_o0 = '1') else
                   sig_10_o0(11);
  sig_13_o0(12) <= sig_16_o0(12) when (sig_14_o0 = '1') else
                   sig_10_o0(12);
  sig_13_o0(13) <= sig_16_o0(13) when (sig_14_o0 = '1') else
                   sig_10_o0(13);
  sig_13_o0(14) <= sig_16_o0(14) when (sig_14_o0 = '1') else
                   sig_10_o0(14);
  sig_13_o0(15) <= sig_16_o0(15) when (sig_14_o0 = '1') else
                   sig_10_o0(15);
  sig_13_o0(16) <= sig_16_o0(16) when (sig_14_o0 = '1') else
                   sig_10_o0(16);
  sig_16_o0(0) <= "" & sig_17_o0;
  sig_16_o0(1) <= "" & sig_93_o0;
  sig_16_o0(2) <= "" & sig_96_o0;
  sig_16_o0(3) <= "" & sig_99_o0;
  sig_16_o0(4) <= "" & sig_102_o0;
  sig_16_o0(5) <= "" & sig_105_o0;
  sig_16_o0(6) <= "" & sig_108_o0;
  sig_16_o0(7) <= "" & sig_111_o0;
  sig_16_o0(8) <= "" & sig_114_o0;
  sig_16_o0(9) <= "" & sig_117_o0;
  sig_16_o0(10) <= "" & sig_120_o0;
  sig_16_o0(11) <= "" & sig_123_o0;
  sig_16_o0(12) <= "" & sig_126_o0;
  sig_16_o0(13) <= "" & sig_129_o0;
  sig_16_o0(14) <= "" & sig_132_o0;
  sig_16_o0(15) <= "" & sig_135_o0;
  sig_16_o0(16) <= "" & sig_138_o0;
  sig_138_o0 <= sig_88_o0 when (sig_139_o0 = '1') else
                sig_140_o0;
  proc446 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_140_o0 <= sig_141_o0;
      end if;
    end if;
  end process proc446;
  sig_141_o0 <= lava_to_std_logic(sig_11_o0(16));
  sig_139_o0 <= lava_to_std_logic(sig_19_o0(16));
  sig_135_o0 <= sig_80_o0 when (sig_78_o0 = '1') else
                sig_136_o0;
  proc450 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_136_o0 <= sig_137_o0;
      end if;
    end if;
  end process proc450;
  sig_137_o0 <= lava_to_std_logic(sig_11_o0(15));
  sig_132_o0 <= sig_76_o0 when (sig_74_o0 = '1') else
                sig_133_o0;
  proc453 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_133_o0 <= sig_134_o0;
      end if;
    end if;
  end process proc453;
  sig_134_o0 <= lava_to_std_logic(sig_11_o0(14));
  sig_129_o0 <= sig_72_o0 when (sig_70_o0 = '1') else
                sig_130_o0;
  proc456 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_130_o0 <= sig_131_o0;
      end if;
    end if;
  end process proc456;
  sig_131_o0 <= lava_to_std_logic(sig_11_o0(13));
  sig_126_o0 <= sig_68_o0 when (sig_66_o0 = '1') else
                sig_127_o0;
  proc459 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_127_o0 <= sig_128_o0;
      end if;
    end if;
  end process proc459;
  sig_128_o0 <= lava_to_std_logic(sig_11_o0(12));
  sig_123_o0 <= sig_64_o0 when (sig_62_o0 = '1') else
                sig_124_o0;
  proc462 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_124_o0 <= sig_125_o0;
      end if;
    end if;
  end process proc462;
  sig_125_o0 <= lava_to_std_logic(sig_11_o0(11));
  sig_120_o0 <= sig_60_o0 when (sig_58_o0 = '1') else
                sig_121_o0;
  proc465 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_121_o0 <= sig_122_o0;
      end if;
    end if;
  end process proc465;
  sig_122_o0 <= lava_to_std_logic(sig_11_o0(10));
  sig_117_o0 <= sig_56_o0 when (sig_54_o0 = '1') else
                sig_118_o0;
  proc468 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_118_o0 <= sig_119_o0;
      end if;
    end if;
  end process proc468;
  sig_119_o0 <= lava_to_std_logic(sig_11_o0(9));
  sig_114_o0 <= sig_52_o0 when (sig_50_o0 = '1') else
                sig_115_o0;
  proc471 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_115_o0 <= sig_116_o0;
      end if;
    end if;
  end process proc471;
  sig_116_o0 <= lava_to_std_logic(sig_11_o0(8));
  sig_111_o0 <= sig_48_o0 when (sig_46_o0 = '1') else
                sig_112_o0;
  proc474 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_112_o0 <= sig_113_o0;
      end if;
    end if;
  end process proc474;
  sig_113_o0 <= lava_to_std_logic(sig_11_o0(7));
  sig_108_o0 <= sig_44_o0 when (sig_42_o0 = '1') else
                sig_109_o0;
  proc477 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_109_o0 <= sig_110_o0;
      end if;
    end if;
  end process proc477;
  sig_110_o0 <= lava_to_std_logic(sig_11_o0(6));
  sig_105_o0 <= sig_40_o0 when (sig_38_o0 = '1') else
                sig_106_o0;
  proc480 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_106_o0 <= sig_107_o0;
      end if;
    end if;
  end process proc480;
  sig_107_o0 <= lava_to_std_logic(sig_11_o0(5));
  sig_102_o0 <= sig_36_o0 when (sig_34_o0 = '1') else
                sig_103_o0;
  proc483 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_103_o0 <= sig_104_o0;
      end if;
    end if;
  end process proc483;
  sig_104_o0 <= lava_to_std_logic(sig_11_o0(4));
  sig_99_o0 <= sig_32_o0 when (sig_30_o0 = '1') else
               sig_100_o0;
  proc486 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_100_o0 <= sig_101_o0;
      end if;
    end if;
  end process proc486;
  sig_101_o0 <= lava_to_std_logic(sig_11_o0(3));
  sig_96_o0 <= sig_28_o0 when (sig_26_o0 = '1') else
               sig_97_o0;
  proc489 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_97_o0 <= sig_98_o0;
      end if;
    end if;
  end process proc489;
  sig_98_o0 <= lava_to_std_logic(sig_11_o0(2));
  sig_93_o0 <= sig_24_o0 when (sig_22_o0 = '1') else
               sig_94_o0;
  proc492 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_94_o0 <= sig_95_o0;
      end if;
    end if;
  end process proc492;
  sig_95_o0 <= lava_to_std_logic(sig_11_o0(1));
  sig_17_o0 <= sig_92_o0 when (sig_18_o0 = '1') else
               sig_90_o0;
  sig_92_o0 <= sig_83_o0(16);
  proc496 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_90_o0 <= sig_91_o0;
      end if;
    end if;
  end process proc496;
  sig_91_o0 <= lava_to_std_logic(sig_11_o0(0));
  sig_18_o0 <= lava_to_std_logic(sig_19_o0(0));
  sig_19_o0(0) <= sig_89_o0(0) when (sig_12_o0 = '1') else
                  sig_20_o0(0);
  sig_19_o0(1) <= sig_89_o0(1) when (sig_12_o0 = '1') else
                  sig_20_o0(1);
  sig_19_o0(2) <= sig_89_o0(2) when (sig_12_o0 = '1') else
                  sig_20_o0(2);
  sig_19_o0(3) <= sig_89_o0(3) when (sig_12_o0 = '1') else
                  sig_20_o0(3);
  sig_19_o0(4) <= sig_89_o0(4) when (sig_12_o0 = '1') else
                  sig_20_o0(4);
  sig_19_o0(5) <= sig_89_o0(5) when (sig_12_o0 = '1') else
                  sig_20_o0(5);
  sig_19_o0(6) <= sig_89_o0(6) when (sig_12_o0 = '1') else
                  sig_20_o0(6);
  sig_19_o0(7) <= sig_89_o0(7) when (sig_12_o0 = '1') else
                  sig_20_o0(7);
  sig_19_o0(8) <= sig_89_o0(8) when (sig_12_o0 = '1') else
                  sig_20_o0(8);
  sig_19_o0(9) <= sig_89_o0(9) when (sig_12_o0 = '1') else
                  sig_20_o0(9);
  sig_19_o0(10) <= sig_89_o0(10) when (sig_12_o0 = '1') else
                   sig_20_o0(10);
  sig_19_o0(11) <= sig_89_o0(11) when (sig_12_o0 = '1') else
                   sig_20_o0(11);
  sig_19_o0(12) <= sig_89_o0(12) when (sig_12_o0 = '1') else
                   sig_20_o0(12);
  sig_19_o0(13) <= sig_89_o0(13) when (sig_12_o0 = '1') else
                   sig_20_o0(13);
  sig_19_o0(14) <= sig_89_o0(14) when (sig_12_o0 = '1') else
                   sig_20_o0(14);
  sig_19_o0(15) <= sig_89_o0(15) when (sig_12_o0 = '1') else
                   sig_20_o0(15);
  sig_19_o0(16) <= sig_89_o0(16) when (sig_12_o0 = '1') else
                   sig_20_o0(16);
  sig_89_o0(0) <= "" & '1';
  sig_89_o0(1) <= "" & '1';
  sig_89_o0(2) <= "" & '1';
  sig_89_o0(3) <= "" & '1';
  sig_89_o0(4) <= "" & '1';
  sig_89_o0(5) <= "" & '1';
  sig_89_o0(6) <= "" & '1';
  sig_89_o0(7) <= "" & '1';
  sig_89_o0(8) <= "" & '1';
  sig_89_o0(9) <= "" & '1';
  sig_89_o0(10) <= "" & '1';
  sig_89_o0(11) <= "" & '1';
  sig_89_o0(12) <= "" & '1';
  sig_89_o0(13) <= "" & '1';
  sig_89_o0(14) <= "" & '1';
  sig_89_o0(15) <= "" & '1';
  sig_89_o0(16) <= "" & '1';
  sig_20_o0(0) <= "" & sig_21_o0;
  sig_20_o0(1) <= "" & sig_25_o0;
  sig_20_o0(2) <= "" & sig_29_o0;
  sig_20_o0(3) <= "" & sig_33_o0;
  sig_20_o0(4) <= "" & sig_37_o0;
  sig_20_o0(5) <= "" & sig_41_o0;
  sig_20_o0(6) <= "" & sig_45_o0;
  sig_20_o0(7) <= "" & sig_49_o0;
  sig_20_o0(8) <= "" & sig_53_o0;
  sig_20_o0(9) <= "" & sig_57_o0;
  sig_20_o0(10) <= "" & sig_61_o0;
  sig_20_o0(11) <= "" & sig_65_o0;
  sig_20_o0(12) <= "" & sig_69_o0;
  sig_20_o0(13) <= "" & sig_73_o0;
  sig_20_o0(14) <= "" & sig_77_o0;
  sig_20_o0(15) <= "" & sig_81_o0;
  sig_20_o0(16) <= "" & sig_81_o0;
  sig_81_o0 <= (sig_82_o0 or sig_87_o0);
  sig_87_o0 <= not(sig_88_o0);
  sig_88_o0 <= lava_to_std_logic(sig_10_o0(15));
  sig_82_o0 <= sig_83_o0(17);
  -- [("i0",16U,(84).o0),("i1",B,(85).o0),("i2",B,(86).o0)];
  sig_83_o0 <= sig_86_o0 & sig_85_o0 & sig_84_o0;
  sig_86_o0 <= out_ready;
  sig_85_o0 <= in_valid;
  sig_84_o0 <= in_x;
  sig_77_o0 <= (sig_78_o0 or sig_79_o0);
  sig_79_o0 <= not(sig_80_o0);
  sig_80_o0 <= lava_to_std_logic(sig_10_o0(14));
  sig_78_o0 <= lava_to_std_logic(sig_19_o0(15));
  sig_73_o0 <= (sig_74_o0 or sig_75_o0);
  sig_75_o0 <= not(sig_76_o0);
  sig_76_o0 <= lava_to_std_logic(sig_10_o0(13));
  sig_74_o0 <= lava_to_std_logic(sig_19_o0(14));
  sig_69_o0 <= (sig_70_o0 or sig_71_o0);
  sig_71_o0 <= not(sig_72_o0);
  sig_72_o0 <= lava_to_std_logic(sig_10_o0(12));
  sig_70_o0 <= lava_to_std_logic(sig_19_o0(13));
  sig_65_o0 <= (sig_66_o0 or sig_67_o0);
  sig_67_o0 <= not(sig_68_o0);
  sig_68_o0 <= lava_to_std_logic(sig_10_o0(11));
  sig_66_o0 <= lava_to_std_logic(sig_19_o0(12));
  sig_61_o0 <= (sig_62_o0 or sig_63_o0);
  sig_63_o0 <= not(sig_64_o0);
  sig_64_o0 <= lava_to_std_logic(sig_10_o0(10));
  sig_62_o0 <= lava_to_std_logic(sig_19_o0(11));
  sig_57_o0 <= (sig_58_o0 or sig_59_o0);
  sig_59_o0 <= not(sig_60_o0);
  sig_60_o0 <= lava_to_std_logic(sig_10_o0(9));
  sig_58_o0 <= lava_to_std_logic(sig_19_o0(10));
  sig_53_o0 <= (sig_54_o0 or sig_55_o0);
  sig_55_o0 <= not(sig_56_o0);
  sig_56_o0 <= lava_to_std_logic(sig_10_o0(8));
  sig_54_o0 <= lava_to_std_logic(sig_19_o0(9));
  sig_49_o0 <= (sig_50_o0 or sig_51_o0);
  sig_51_o0 <= not(sig_52_o0);
  sig_52_o0 <= lava_to_std_logic(sig_10_o0(7));
  sig_50_o0 <= lava_to_std_logic(sig_19_o0(8));
  sig_45_o0 <= (sig_46_o0 or sig_47_o0);
  sig_47_o0 <= not(sig_48_o0);
  sig_48_o0 <= lava_to_std_logic(sig_10_o0(6));
  sig_46_o0 <= lava_to_std_logic(sig_19_o0(7));
  sig_41_o0 <= (sig_42_o0 or sig_43_o0);
  sig_43_o0 <= not(sig_44_o0);
  sig_44_o0 <= lava_to_std_logic(sig_10_o0(5));
  sig_42_o0 <= lava_to_std_logic(sig_19_o0(6));
  sig_37_o0 <= (sig_38_o0 or sig_39_o0);
  sig_39_o0 <= not(sig_40_o0);
  sig_40_o0 <= lava_to_std_logic(sig_10_o0(4));
  sig_38_o0 <= lava_to_std_logic(sig_19_o0(5));
  sig_33_o0 <= (sig_34_o0 or sig_35_o0);
  sig_35_o0 <= not(sig_36_o0);
  sig_36_o0 <= lava_to_std_logic(sig_10_o0(3));
  sig_34_o0 <= lava_to_std_logic(sig_19_o0(4));
  sig_29_o0 <= (sig_30_o0 or sig_31_o0);
  sig_31_o0 <= not(sig_32_o0);
  sig_32_o0 <= lava_to_std_logic(sig_10_o0(2));
  sig_30_o0 <= lava_to_std_logic(sig_19_o0(3));
  sig_25_o0 <= (sig_26_o0 or sig_27_o0);
  sig_27_o0 <= not(sig_28_o0);
  sig_28_o0 <= lava_to_std_logic(sig_10_o0(1));
  sig_26_o0 <= lava_to_std_logic(sig_19_o0(2));
  sig_21_o0 <= (sig_22_o0 or sig_23_o0);
  sig_23_o0 <= not(sig_24_o0);
  sig_24_o0 <= lava_to_std_logic(sig_10_o0(0));
  sig_22_o0 <= lava_to_std_logic(sig_19_o0(1));
  sig_14_o0 <= not(sig_15_o0);
  sig_15_o0 <= (sig_12_o0 or '0');
  sig_12_o0 <= reset;
  out_valid <= sig_2_o0;
  in_ready <= sig_235_o0;
  out_x <= sig_237_o0;
end architecture str;
