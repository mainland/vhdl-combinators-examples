library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.lava.all;
use work.all;
entity incrementer is
  port(clk : in std_logic;
       in_x : in std_logic_vector(15 downto 0);
       reset : in std_logic;
       in_valid : in std_logic;
       out_ready : in std_logic;
       out_valid : out std_logic;
       in_ready : out std_logic;
       out_x : out std_logic_vector(15 downto 0));
end entity incrementer;
architecture str of incrementer is
  signal sig_271_o0 : std_logic_vector(15 downto 0);
  signal sig_272_o0 : std_logic_vector(15 downto 0);
  signal sig_269_o0 : std_logic;
  signal sig_270_o0 : std_logic;
  signal sig_2_o0 : std_logic;
  signal sig_3_o0 : std_logic;
  signal sig_4_o0 : std_logic_vector(17 downto 0);
  signal sig_268_o0 : std_logic;
  signal sig_5_o0 : std_logic_vector(15 downto 0);
  signal sig_6_o0 : std_logic_vector(16 downto 0);
  signal sig_267_o0 : std_logic_vector(15 downto 0);
  signal sig_7_o0 : std_logic;
  signal sig_8_o0 : std_logic_vector(16 downto 0);
  signal sig_170_o0 : std_logic_vector(15 downto 0);
  signal sig_174_o0 : std_logic_vector(15 downto 0);
  signal sig_175_o0 : std_logic_vector(15 downto 0);
  signal sig_176_o0 : std_logic_vector(15 downto 0);
  signal sig_180_o0 : std_logic_vector(15 downto 0);
  signal sig_181_o0 : std_logic_vector(15 downto 0);
  signal sig_182_o0 : std_logic_vector(15 downto 0);
  signal sig_186_o0 : std_logic_vector(15 downto 0);
  signal sig_187_o0 : std_logic_vector(15 downto 0);
  signal sig_188_o0 : std_logic_vector(15 downto 0);
  signal sig_192_o0 : std_logic_vector(15 downto 0);
  signal sig_193_o0 : std_logic_vector(15 downto 0);
  signal sig_194_o0 : std_logic_vector(15 downto 0);
  signal sig_198_o0 : std_logic_vector(15 downto 0);
  signal sig_199_o0 : std_logic_vector(15 downto 0);
  signal sig_200_o0 : std_logic_vector(15 downto 0);
  signal sig_204_o0 : std_logic_vector(15 downto 0);
  signal sig_205_o0 : std_logic_vector(15 downto 0);
  signal sig_206_o0 : std_logic_vector(15 downto 0);
  signal sig_210_o0 : std_logic_vector(15 downto 0);
  signal sig_211_o0 : std_logic_vector(15 downto 0);
  signal sig_212_o0 : std_logic_vector(15 downto 0);
  signal sig_216_o0 : std_logic_vector(15 downto 0);
  signal sig_217_o0 : std_logic_vector(15 downto 0);
  signal sig_218_o0 : std_logic_vector(15 downto 0);
  signal sig_222_o0 : std_logic_vector(15 downto 0);
  signal sig_223_o0 : std_logic_vector(15 downto 0);
  signal sig_224_o0 : std_logic_vector(15 downto 0);
  signal sig_228_o0 : std_logic_vector(15 downto 0);
  signal sig_229_o0 : std_logic_vector(15 downto 0);
  signal sig_230_o0 : std_logic_vector(15 downto 0);
  signal sig_234_o0 : std_logic_vector(15 downto 0);
  signal sig_235_o0 : std_logic_vector(15 downto 0);
  signal sig_236_o0 : std_logic_vector(15 downto 0);
  signal sig_240_o0 : std_logic_vector(15 downto 0);
  signal sig_241_o0 : std_logic_vector(15 downto 0);
  signal sig_242_o0 : std_logic_vector(15 downto 0);
  signal sig_246_o0 : std_logic_vector(15 downto 0);
  signal sig_247_o0 : std_logic_vector(15 downto 0);
  signal sig_248_o0 : std_logic_vector(15 downto 0);
  signal sig_252_o0 : std_logic_vector(15 downto 0);
  signal sig_253_o0 : std_logic_vector(15 downto 0);
  signal sig_254_o0 : std_logic_vector(15 downto 0);
  signal sig_258_o0 : std_logic_vector(15 downto 0);
  signal sig_259_o0 : std_logic_vector(15 downto 0);
  signal sig_260_o0 : std_logic_vector(15 downto 0);
  signal sig_264_o0 : std_logic_vector(15 downto 0);
  signal sig_265_o0 : std_logic_vector(15 downto 0);
  signal sig_266_o0 : std_logic_vector(15 downto 0);
  signal sig_263_o0 : std_logic_vector(15 downto 0);
  signal sig_261_o0 : std_logic;
  signal sig_262_o0 : std_logic;
  signal sig_257_o0 : std_logic_vector(15 downto 0);
  signal sig_255_o0 : std_logic;
  signal sig_256_o0 : std_logic;
  signal sig_251_o0 : std_logic_vector(15 downto 0);
  signal sig_249_o0 : std_logic;
  signal sig_250_o0 : std_logic;
  signal sig_245_o0 : std_logic_vector(15 downto 0);
  signal sig_243_o0 : std_logic;
  signal sig_244_o0 : std_logic;
  signal sig_239_o0 : std_logic_vector(15 downto 0);
  signal sig_237_o0 : std_logic;
  signal sig_238_o0 : std_logic;
  signal sig_233_o0 : std_logic_vector(15 downto 0);
  signal sig_231_o0 : std_logic;
  signal sig_232_o0 : std_logic;
  signal sig_227_o0 : std_logic_vector(15 downto 0);
  signal sig_225_o0 : std_logic;
  signal sig_226_o0 : std_logic;
  signal sig_221_o0 : std_logic_vector(15 downto 0);
  signal sig_219_o0 : std_logic;
  signal sig_220_o0 : std_logic;
  signal sig_215_o0 : std_logic_vector(15 downto 0);
  signal sig_213_o0 : std_logic;
  signal sig_214_o0 : std_logic;
  signal sig_209_o0 : std_logic_vector(15 downto 0);
  signal sig_207_o0 : std_logic;
  signal sig_208_o0 : std_logic;
  signal sig_203_o0 : std_logic_vector(15 downto 0);
  signal sig_201_o0 : std_logic;
  signal sig_202_o0 : std_logic;
  signal sig_197_o0 : std_logic_vector(15 downto 0);
  signal sig_195_o0 : std_logic;
  signal sig_196_o0 : std_logic;
  signal sig_191_o0 : std_logic_vector(15 downto 0);
  signal sig_189_o0 : std_logic;
  signal sig_190_o0 : std_logic;
  signal sig_185_o0 : std_logic_vector(15 downto 0);
  signal sig_183_o0 : std_logic;
  signal sig_184_o0 : std_logic;
  signal sig_179_o0 : std_logic_vector(15 downto 0);
  signal sig_177_o0 : std_logic;
  signal sig_178_o0 : std_logic;
  signal sig_173_o0 : std_logic_vector(15 downto 0);
  signal sig_171_o0 : std_logic;
  signal sig_172_o0 : std_logic;
  signal sig_9_o0 : std_logic;
  signal sig_11_o0 : std_logic;
  signal sig_33_o0 : std_logic;
  signal sig_34_o0 : std_logic;
  signal sig_42_o0 : std_logic;
  signal sig_43_o0 : std_logic;
  signal sig_51_o0 : std_logic;
  signal sig_52_o0 : std_logic;
  signal sig_60_o0 : std_logic;
  signal sig_61_o0 : std_logic;
  signal sig_69_o0 : std_logic;
  signal sig_70_o0 : std_logic;
  signal sig_78_o0 : std_logic;
  signal sig_79_o0 : std_logic;
  signal sig_87_o0 : std_logic;
  signal sig_88_o0 : std_logic;
  signal sig_96_o0 : std_logic;
  signal sig_97_o0 : std_logic;
  signal sig_105_o0 : std_logic;
  signal sig_106_o0 : std_logic;
  signal sig_114_o0 : std_logic;
  signal sig_115_o0 : std_logic;
  signal sig_123_o0 : std_logic;
  signal sig_124_o0 : std_logic;
  signal sig_132_o0 : std_logic;
  signal sig_133_o0 : std_logic;
  signal sig_141_o0 : std_logic;
  signal sig_142_o0 : std_logic;
  signal sig_150_o0 : std_logic;
  signal sig_151_o0 : std_logic;
  signal sig_159_o0 : std_logic;
  signal sig_160_o0 : std_logic;
  signal sig_168_o0 : std_logic;
  signal sig_169_o0 : std_logic;
  signal sig_167_o0 : std_logic;
  signal sig_161_o0 : std_logic;
  signal sig_162_o0 : std_logic;
  signal sig_163_o0 : std_logic;
  signal sig_164_o0 : std_logic;
  signal sig_165_o0 : std_logic;
  signal sig_166_o0 : std_logic;
  signal sig_158_o0 : std_logic;
  signal sig_152_o0 : std_logic;
  signal sig_153_o0 : std_logic;
  signal sig_154_o0 : std_logic;
  signal sig_155_o0 : std_logic;
  signal sig_156_o0 : std_logic;
  signal sig_157_o0 : std_logic;
  signal sig_149_o0 : std_logic;
  signal sig_143_o0 : std_logic;
  signal sig_144_o0 : std_logic;
  signal sig_145_o0 : std_logic;
  signal sig_146_o0 : std_logic;
  signal sig_147_o0 : std_logic;
  signal sig_148_o0 : std_logic;
  signal sig_140_o0 : std_logic;
  signal sig_134_o0 : std_logic;
  signal sig_135_o0 : std_logic;
  signal sig_136_o0 : std_logic;
  signal sig_137_o0 : std_logic;
  signal sig_138_o0 : std_logic;
  signal sig_139_o0 : std_logic;
  signal sig_131_o0 : std_logic;
  signal sig_125_o0 : std_logic;
  signal sig_126_o0 : std_logic;
  signal sig_127_o0 : std_logic;
  signal sig_128_o0 : std_logic;
  signal sig_129_o0 : std_logic;
  signal sig_130_o0 : std_logic;
  signal sig_122_o0 : std_logic;
  signal sig_116_o0 : std_logic;
  signal sig_117_o0 : std_logic;
  signal sig_118_o0 : std_logic;
  signal sig_119_o0 : std_logic;
  signal sig_120_o0 : std_logic;
  signal sig_121_o0 : std_logic;
  signal sig_113_o0 : std_logic;
  signal sig_107_o0 : std_logic;
  signal sig_108_o0 : std_logic;
  signal sig_109_o0 : std_logic;
  signal sig_110_o0 : std_logic;
  signal sig_111_o0 : std_logic;
  signal sig_112_o0 : std_logic;
  signal sig_104_o0 : std_logic;
  signal sig_98_o0 : std_logic;
  signal sig_99_o0 : std_logic;
  signal sig_100_o0 : std_logic;
  signal sig_101_o0 : std_logic;
  signal sig_102_o0 : std_logic;
  signal sig_103_o0 : std_logic;
  signal sig_95_o0 : std_logic;
  signal sig_89_o0 : std_logic;
  signal sig_90_o0 : std_logic;
  signal sig_91_o0 : std_logic;
  signal sig_92_o0 : std_logic;
  signal sig_93_o0 : std_logic;
  signal sig_94_o0 : std_logic;
  signal sig_86_o0 : std_logic;
  signal sig_80_o0 : std_logic;
  signal sig_81_o0 : std_logic;
  signal sig_82_o0 : std_logic;
  signal sig_83_o0 : std_logic;
  signal sig_84_o0 : std_logic;
  signal sig_85_o0 : std_logic;
  signal sig_77_o0 : std_logic;
  signal sig_71_o0 : std_logic;
  signal sig_72_o0 : std_logic;
  signal sig_73_o0 : std_logic;
  signal sig_74_o0 : std_logic;
  signal sig_75_o0 : std_logic;
  signal sig_76_o0 : std_logic;
  signal sig_68_o0 : std_logic;
  signal sig_62_o0 : std_logic;
  signal sig_63_o0 : std_logic;
  signal sig_64_o0 : std_logic;
  signal sig_65_o0 : std_logic;
  signal sig_66_o0 : std_logic;
  signal sig_67_o0 : std_logic;
  signal sig_59_o0 : std_logic;
  signal sig_53_o0 : std_logic;
  signal sig_54_o0 : std_logic;
  signal sig_55_o0 : std_logic;
  signal sig_56_o0 : std_logic;
  signal sig_57_o0 : std_logic;
  signal sig_58_o0 : std_logic;
  signal sig_50_o0 : std_logic;
  signal sig_44_o0 : std_logic;
  signal sig_45_o0 : std_logic;
  signal sig_46_o0 : std_logic;
  signal sig_47_o0 : std_logic;
  signal sig_48_o0 : std_logic;
  signal sig_49_o0 : std_logic;
  signal sig_41_o0 : std_logic;
  signal sig_35_o0 : std_logic;
  signal sig_36_o0 : std_logic;
  signal sig_37_o0 : std_logic;
  signal sig_38_o0 : std_logic;
  signal sig_39_o0 : std_logic;
  signal sig_40_o0 : std_logic;
  signal sig_32_o0 : std_logic;
  signal sig_12_o0 : std_logic;
  signal sig_14_o0 : std_logic;
  signal sig_15_o0 : std_logic;
  signal sig_16_o0 : std_logic;
  signal sig_31_o0 : std_logic;
  signal sig_17_o0 : std_logic;
  signal sig_23_o0 : std_logic;
  signal sig_24_o0 : std_logic;
  signal sig_25_o0 : std_logic;
  signal sig_30_o0 : std_logic;
  signal sig_29_o0 : std_logic;
  signal sig_26_o0 : std_logic;
  signal sig_27_o0 : std_logic;
  signal sig_28_o0 : std_logic;
  signal sig_18_o0 : std_logic;
  signal sig_19_o0 : std_logic_vector(17 downto 0);
  signal sig_22_o0 : std_logic;
  signal sig_21_o0 : std_logic;
  signal sig_20_o0 : std_logic_vector(15 downto 0);
  signal sig_13_o0 : std_logic;
  signal sig_10_o0 : std_logic;
begin
  sig_271_o0 <= sig_272_o0;
  sig_272_o0 <= sig_4_o0(15 downto 0);
  sig_269_o0 <= sig_270_o0;
  sig_270_o0 <= sig_4_o0(17);
  sig_2_o0 <= sig_3_o0;
  sig_3_o0 <= sig_4_o0(16);
  -- [("i0",16U,(5).o0),("i1",B,(268).o0),("i2",B,(163).o0)];
  sig_4_o0 <= sig_163_o0 & sig_268_o0 & sig_5_o0;
  sig_268_o0 <= sig_6_o0(0);
  sig_5_o0 <= sig_6_o0(16 downto 1);
  -- [("i0",B,(7).o0),("i1",16U,(267).o0)];
  sig_6_o0 <= sig_267_o0 & sig_7_o0;
  sig_267_o0 <= sig_8_o0(16 downto 1);
  sig_7_o0 <= sig_8_o0(0);
  -- [("i0",B,(9).o0),("i1",16U,(170).o0)];
  sig_8_o0 <= sig_170_o0 & sig_9_o0;
  sig_170_o0 <= sig_174_o0 when (sig_171_o0 = '1') else
                sig_173_o0;
  sig_174_o0 <= std_logic_vector((unsigned(sig_175_o0) + to_unsigned(1,
                                                                     16)));
  proc289 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_175_o0 <= sig_176_o0;
      end if;
    end if;
  end process proc289;
  sig_176_o0 <= sig_180_o0 when (sig_177_o0 = '1') else
                sig_179_o0;
  sig_180_o0 <= std_logic_vector((unsigned(sig_181_o0) + to_unsigned(1,
                                                                     16)));
  proc292 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_181_o0 <= sig_182_o0;
      end if;
    end if;
  end process proc292;
  sig_182_o0 <= sig_186_o0 when (sig_183_o0 = '1') else
                sig_185_o0;
  sig_186_o0 <= std_logic_vector((unsigned(sig_187_o0) + to_unsigned(1,
                                                                     16)));
  proc295 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_187_o0 <= sig_188_o0;
      end if;
    end if;
  end process proc295;
  sig_188_o0 <= sig_192_o0 when (sig_189_o0 = '1') else
                sig_191_o0;
  sig_192_o0 <= std_logic_vector((unsigned(sig_193_o0) + to_unsigned(1,
                                                                     16)));
  proc298 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_193_o0 <= sig_194_o0;
      end if;
    end if;
  end process proc298;
  sig_194_o0 <= sig_198_o0 when (sig_195_o0 = '1') else
                sig_197_o0;
  sig_198_o0 <= std_logic_vector((unsigned(sig_199_o0) + to_unsigned(1,
                                                                     16)));
  proc301 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_199_o0 <= sig_200_o0;
      end if;
    end if;
  end process proc301;
  sig_200_o0 <= sig_204_o0 when (sig_201_o0 = '1') else
                sig_203_o0;
  sig_204_o0 <= std_logic_vector((unsigned(sig_205_o0) + to_unsigned(1,
                                                                     16)));
  proc304 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_205_o0 <= sig_206_o0;
      end if;
    end if;
  end process proc304;
  sig_206_o0 <= sig_210_o0 when (sig_207_o0 = '1') else
                sig_209_o0;
  sig_210_o0 <= std_logic_vector((unsigned(sig_211_o0) + to_unsigned(1,
                                                                     16)));
  proc307 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_211_o0 <= sig_212_o0;
      end if;
    end if;
  end process proc307;
  sig_212_o0 <= sig_216_o0 when (sig_213_o0 = '1') else
                sig_215_o0;
  sig_216_o0 <= std_logic_vector((unsigned(sig_217_o0) + to_unsigned(1,
                                                                     16)));
  proc310 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_217_o0 <= sig_218_o0;
      end if;
    end if;
  end process proc310;
  sig_218_o0 <= sig_222_o0 when (sig_219_o0 = '1') else
                sig_221_o0;
  sig_222_o0 <= std_logic_vector((unsigned(sig_223_o0) + to_unsigned(1,
                                                                     16)));
  proc313 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_223_o0 <= sig_224_o0;
      end if;
    end if;
  end process proc313;
  sig_224_o0 <= sig_228_o0 when (sig_225_o0 = '1') else
                sig_227_o0;
  sig_228_o0 <= std_logic_vector((unsigned(sig_229_o0) + to_unsigned(1,
                                                                     16)));
  proc316 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_229_o0 <= sig_230_o0;
      end if;
    end if;
  end process proc316;
  sig_230_o0 <= sig_234_o0 when (sig_231_o0 = '1') else
                sig_233_o0;
  sig_234_o0 <= std_logic_vector((unsigned(sig_235_o0) + to_unsigned(1,
                                                                     16)));
  proc319 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_235_o0 <= sig_236_o0;
      end if;
    end if;
  end process proc319;
  sig_236_o0 <= sig_240_o0 when (sig_237_o0 = '1') else
                sig_239_o0;
  sig_240_o0 <= std_logic_vector((unsigned(sig_241_o0) + to_unsigned(1,
                                                                     16)));
  proc322 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_241_o0 <= sig_242_o0;
      end if;
    end if;
  end process proc322;
  sig_242_o0 <= sig_246_o0 when (sig_243_o0 = '1') else
                sig_245_o0;
  sig_246_o0 <= std_logic_vector((unsigned(sig_247_o0) + to_unsigned(1,
                                                                     16)));
  proc325 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_247_o0 <= sig_248_o0;
      end if;
    end if;
  end process proc325;
  sig_248_o0 <= sig_252_o0 when (sig_249_o0 = '1') else
                sig_251_o0;
  sig_252_o0 <= std_logic_vector((unsigned(sig_253_o0) + to_unsigned(1,
                                                                     16)));
  proc328 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_253_o0 <= sig_254_o0;
      end if;
    end if;
  end process proc328;
  sig_254_o0 <= sig_258_o0 when (sig_255_o0 = '1') else
                sig_257_o0;
  sig_258_o0 <= std_logic_vector((unsigned(sig_259_o0) + to_unsigned(1,
                                                                     16)));
  proc331 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_259_o0 <= sig_260_o0;
      end if;
    end if;
  end process proc331;
  sig_260_o0 <= sig_264_o0 when (sig_261_o0 = '1') else
                sig_263_o0;
  sig_264_o0 <= std_logic_vector((unsigned(sig_265_o0) + to_unsigned(1,
                                                                     16)));
  proc334 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_265_o0 <= sig_266_o0;
      end if;
    end if;
  end process proc334;
  sig_266_o0 <= sig_19_o0(15 downto 0);
  proc336 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_263_o0 <= sig_260_o0;
      end if;
    end if;
  end process proc336;
  sig_261_o0 <= (sig_13_o0 and sig_262_o0);
  proc338 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_262_o0 <= sig_163_o0;
      end if;
    end if;
  end process proc338;
  proc339 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_257_o0 <= sig_254_o0;
      end if;
    end if;
  end process proc339;
  sig_255_o0 <= (sig_13_o0 and sig_256_o0);
  proc341 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_256_o0 <= sig_154_o0;
      end if;
    end if;
  end process proc341;
  proc342 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_251_o0 <= sig_248_o0;
      end if;
    end if;
  end process proc342;
  sig_249_o0 <= (sig_13_o0 and sig_250_o0);
  proc344 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_250_o0 <= sig_145_o0;
      end if;
    end if;
  end process proc344;
  proc345 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_245_o0 <= sig_242_o0;
      end if;
    end if;
  end process proc345;
  sig_243_o0 <= (sig_13_o0 and sig_244_o0);
  proc347 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_244_o0 <= sig_136_o0;
      end if;
    end if;
  end process proc347;
  proc348 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_239_o0 <= sig_236_o0;
      end if;
    end if;
  end process proc348;
  sig_237_o0 <= (sig_13_o0 and sig_238_o0);
  proc350 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_238_o0 <= sig_127_o0;
      end if;
    end if;
  end process proc350;
  proc351 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_233_o0 <= sig_230_o0;
      end if;
    end if;
  end process proc351;
  sig_231_o0 <= (sig_13_o0 and sig_232_o0);
  proc353 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_232_o0 <= sig_118_o0;
      end if;
    end if;
  end process proc353;
  proc354 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_227_o0 <= sig_224_o0;
      end if;
    end if;
  end process proc354;
  sig_225_o0 <= (sig_13_o0 and sig_226_o0);
  proc356 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_226_o0 <= sig_109_o0;
      end if;
    end if;
  end process proc356;
  proc357 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_221_o0 <= sig_218_o0;
      end if;
    end if;
  end process proc357;
  sig_219_o0 <= (sig_13_o0 and sig_220_o0);
  proc359 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_220_o0 <= sig_100_o0;
      end if;
    end if;
  end process proc359;
  proc360 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_215_o0 <= sig_212_o0;
      end if;
    end if;
  end process proc360;
  sig_213_o0 <= (sig_13_o0 and sig_214_o0);
  proc362 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_214_o0 <= sig_91_o0;
      end if;
    end if;
  end process proc362;
  proc363 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_209_o0 <= sig_206_o0;
      end if;
    end if;
  end process proc363;
  sig_207_o0 <= (sig_13_o0 and sig_208_o0);
  proc365 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_208_o0 <= sig_82_o0;
      end if;
    end if;
  end process proc365;
  proc366 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_203_o0 <= sig_200_o0;
      end if;
    end if;
  end process proc366;
  sig_201_o0 <= (sig_13_o0 and sig_202_o0);
  proc368 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_202_o0 <= sig_73_o0;
      end if;
    end if;
  end process proc368;
  proc369 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_197_o0 <= sig_194_o0;
      end if;
    end if;
  end process proc369;
  sig_195_o0 <= (sig_13_o0 and sig_196_o0);
  proc371 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_196_o0 <= sig_64_o0;
      end if;
    end if;
  end process proc371;
  proc372 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_191_o0 <= sig_188_o0;
      end if;
    end if;
  end process proc372;
  sig_189_o0 <= (sig_13_o0 and sig_190_o0);
  proc374 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_190_o0 <= sig_55_o0;
      end if;
    end if;
  end process proc374;
  proc375 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_185_o0 <= sig_182_o0;
      end if;
    end if;
  end process proc375;
  sig_183_o0 <= (sig_13_o0 and sig_184_o0);
  proc377 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_184_o0 <= sig_46_o0;
      end if;
    end if;
  end process proc377;
  proc378 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_179_o0 <= sig_176_o0;
      end if;
    end if;
  end process proc378;
  sig_177_o0 <= (sig_13_o0 and sig_178_o0);
  proc380 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_178_o0 <= sig_37_o0;
      end if;
    end if;
  end process proc380;
  proc381 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_173_o0 <= sig_170_o0;
      end if;
    end if;
  end process proc381;
  sig_171_o0 <= (sig_13_o0 and sig_172_o0);
  proc383 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_172_o0 <= sig_15_o0;
      end if;
    end if;
  end process proc383;
  sig_9_o0 <= '0' when (sig_10_o0 = '1') else
              sig_11_o0;
  sig_11_o0 <= sig_33_o0 when (sig_12_o0 = '1') else
               sig_32_o0;
  proc386 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_33_o0 <= sig_34_o0;
      end if;
    end if;
  end process proc386;
  sig_34_o0 <= sig_42_o0 when (sig_35_o0 = '1') else
               sig_41_o0;
  proc388 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_42_o0 <= sig_43_o0;
      end if;
    end if;
  end process proc388;
  sig_43_o0 <= sig_51_o0 when (sig_44_o0 = '1') else
               sig_50_o0;
  proc390 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_51_o0 <= sig_52_o0;
      end if;
    end if;
  end process proc390;
  sig_52_o0 <= sig_60_o0 when (sig_53_o0 = '1') else
               sig_59_o0;
  proc392 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_60_o0 <= sig_61_o0;
      end if;
    end if;
  end process proc392;
  sig_61_o0 <= sig_69_o0 when (sig_62_o0 = '1') else
               sig_68_o0;
  proc394 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_69_o0 <= sig_70_o0;
      end if;
    end if;
  end process proc394;
  sig_70_o0 <= sig_78_o0 when (sig_71_o0 = '1') else
               sig_77_o0;
  proc396 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_78_o0 <= sig_79_o0;
      end if;
    end if;
  end process proc396;
  sig_79_o0 <= sig_87_o0 when (sig_80_o0 = '1') else
               sig_86_o0;
  proc398 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_87_o0 <= sig_88_o0;
      end if;
    end if;
  end process proc398;
  sig_88_o0 <= sig_96_o0 when (sig_89_o0 = '1') else
               sig_95_o0;
  proc400 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_96_o0 <= sig_97_o0;
      end if;
    end if;
  end process proc400;
  sig_97_o0 <= sig_105_o0 when (sig_98_o0 = '1') else
               sig_104_o0;
  proc402 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_105_o0 <= sig_106_o0;
      end if;
    end if;
  end process proc402;
  sig_106_o0 <= sig_114_o0 when (sig_107_o0 = '1') else
                sig_113_o0;
  proc404 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_114_o0 <= sig_115_o0;
      end if;
    end if;
  end process proc404;
  sig_115_o0 <= sig_123_o0 when (sig_116_o0 = '1') else
                sig_122_o0;
  proc406 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_123_o0 <= sig_124_o0;
      end if;
    end if;
  end process proc406;
  sig_124_o0 <= sig_132_o0 when (sig_125_o0 = '1') else
                sig_131_o0;
  proc408 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_132_o0 <= sig_133_o0;
      end if;
    end if;
  end process proc408;
  sig_133_o0 <= sig_141_o0 when (sig_134_o0 = '1') else
                sig_140_o0;
  proc410 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_141_o0 <= sig_142_o0;
      end if;
    end if;
  end process proc410;
  sig_142_o0 <= sig_150_o0 when (sig_143_o0 = '1') else
                sig_149_o0;
  proc412 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_150_o0 <= sig_151_o0;
      end if;
    end if;
  end process proc412;
  sig_151_o0 <= sig_159_o0 when (sig_152_o0 = '1') else
                sig_158_o0;
  proc414 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_159_o0 <= sig_160_o0;
      end if;
    end if;
  end process proc414;
  sig_160_o0 <= sig_168_o0 when (sig_161_o0 = '1') else
                sig_167_o0;
  proc416 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_168_o0 <= sig_169_o0;
      end if;
    end if;
  end process proc416;
  sig_169_o0 <= sig_19_o0(16);
  proc418 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_167_o0 <= sig_160_o0;
      end if;
    end if;
  end process proc418;
  sig_161_o0 <= (sig_13_o0 and sig_162_o0);
  proc420 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_162_o0 <= sig_163_o0;
      end if;
    end if;
  end process proc420;
  sig_163_o0 <= '1' when (sig_10_o0 = '1') else
                sig_164_o0;
  sig_164_o0 <= (sig_155_o0 or sig_165_o0);
  sig_165_o0 <= not(sig_166_o0);
  sig_166_o0 <= '0' when (sig_10_o0 = '1') else
                sig_160_o0;
  proc425 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_158_o0 <= sig_151_o0;
      end if;
    end if;
  end process proc425;
  sig_152_o0 <= (sig_13_o0 and sig_153_o0);
  proc427 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_153_o0 <= sig_154_o0;
      end if;
    end if;
  end process proc427;
  sig_154_o0 <= '1' when (sig_10_o0 = '1') else
                sig_155_o0;
  sig_155_o0 <= (sig_146_o0 or sig_156_o0);
  sig_156_o0 <= not(sig_157_o0);
  sig_157_o0 <= '0' when (sig_10_o0 = '1') else
                sig_151_o0;
  proc432 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_149_o0 <= sig_142_o0;
      end if;
    end if;
  end process proc432;
  sig_143_o0 <= (sig_13_o0 and sig_144_o0);
  proc434 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_144_o0 <= sig_145_o0;
      end if;
    end if;
  end process proc434;
  sig_145_o0 <= '1' when (sig_10_o0 = '1') else
                sig_146_o0;
  sig_146_o0 <= (sig_137_o0 or sig_147_o0);
  sig_147_o0 <= not(sig_148_o0);
  sig_148_o0 <= '0' when (sig_10_o0 = '1') else
                sig_142_o0;
  proc439 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_140_o0 <= sig_133_o0;
      end if;
    end if;
  end process proc439;
  sig_134_o0 <= (sig_13_o0 and sig_135_o0);
  proc441 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_135_o0 <= sig_136_o0;
      end if;
    end if;
  end process proc441;
  sig_136_o0 <= '1' when (sig_10_o0 = '1') else
                sig_137_o0;
  sig_137_o0 <= (sig_128_o0 or sig_138_o0);
  sig_138_o0 <= not(sig_139_o0);
  sig_139_o0 <= '0' when (sig_10_o0 = '1') else
                sig_133_o0;
  proc446 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_131_o0 <= sig_124_o0;
      end if;
    end if;
  end process proc446;
  sig_125_o0 <= (sig_13_o0 and sig_126_o0);
  proc448 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_126_o0 <= sig_127_o0;
      end if;
    end if;
  end process proc448;
  sig_127_o0 <= '1' when (sig_10_o0 = '1') else
                sig_128_o0;
  sig_128_o0 <= (sig_119_o0 or sig_129_o0);
  sig_129_o0 <= not(sig_130_o0);
  sig_130_o0 <= '0' when (sig_10_o0 = '1') else
                sig_124_o0;
  proc453 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_122_o0 <= sig_115_o0;
      end if;
    end if;
  end process proc453;
  sig_116_o0 <= (sig_13_o0 and sig_117_o0);
  proc455 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_117_o0 <= sig_118_o0;
      end if;
    end if;
  end process proc455;
  sig_118_o0 <= '1' when (sig_10_o0 = '1') else
                sig_119_o0;
  sig_119_o0 <= (sig_110_o0 or sig_120_o0);
  sig_120_o0 <= not(sig_121_o0);
  sig_121_o0 <= '0' when (sig_10_o0 = '1') else
                sig_115_o0;
  proc460 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_113_o0 <= sig_106_o0;
      end if;
    end if;
  end process proc460;
  sig_107_o0 <= (sig_13_o0 and sig_108_o0);
  proc462 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_108_o0 <= sig_109_o0;
      end if;
    end if;
  end process proc462;
  sig_109_o0 <= '1' when (sig_10_o0 = '1') else
                sig_110_o0;
  sig_110_o0 <= (sig_101_o0 or sig_111_o0);
  sig_111_o0 <= not(sig_112_o0);
  sig_112_o0 <= '0' when (sig_10_o0 = '1') else
                sig_106_o0;
  proc467 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_104_o0 <= sig_97_o0;
      end if;
    end if;
  end process proc467;
  sig_98_o0 <= (sig_13_o0 and sig_99_o0);
  proc469 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_99_o0 <= sig_100_o0;
      end if;
    end if;
  end process proc469;
  sig_100_o0 <= '1' when (sig_10_o0 = '1') else
                sig_101_o0;
  sig_101_o0 <= (sig_92_o0 or sig_102_o0);
  sig_102_o0 <= not(sig_103_o0);
  sig_103_o0 <= '0' when (sig_10_o0 = '1') else
                sig_97_o0;
  proc474 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_95_o0 <= sig_88_o0;
      end if;
    end if;
  end process proc474;
  sig_89_o0 <= (sig_13_o0 and sig_90_o0);
  proc476 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_90_o0 <= sig_91_o0;
      end if;
    end if;
  end process proc476;
  sig_91_o0 <= '1' when (sig_10_o0 = '1') else
               sig_92_o0;
  sig_92_o0 <= (sig_83_o0 or sig_93_o0);
  sig_93_o0 <= not(sig_94_o0);
  sig_94_o0 <= '0' when (sig_10_o0 = '1') else
               sig_88_o0;
  proc481 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_86_o0 <= sig_79_o0;
      end if;
    end if;
  end process proc481;
  sig_80_o0 <= (sig_13_o0 and sig_81_o0);
  proc483 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_81_o0 <= sig_82_o0;
      end if;
    end if;
  end process proc483;
  sig_82_o0 <= '1' when (sig_10_o0 = '1') else
               sig_83_o0;
  sig_83_o0 <= (sig_74_o0 or sig_84_o0);
  sig_84_o0 <= not(sig_85_o0);
  sig_85_o0 <= '0' when (sig_10_o0 = '1') else
               sig_79_o0;
  proc488 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_77_o0 <= sig_70_o0;
      end if;
    end if;
  end process proc488;
  sig_71_o0 <= (sig_13_o0 and sig_72_o0);
  proc490 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_72_o0 <= sig_73_o0;
      end if;
    end if;
  end process proc490;
  sig_73_o0 <= '1' when (sig_10_o0 = '1') else
               sig_74_o0;
  sig_74_o0 <= (sig_65_o0 or sig_75_o0);
  sig_75_o0 <= not(sig_76_o0);
  sig_76_o0 <= '0' when (sig_10_o0 = '1') else
               sig_70_o0;
  proc495 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_68_o0 <= sig_61_o0;
      end if;
    end if;
  end process proc495;
  sig_62_o0 <= (sig_13_o0 and sig_63_o0);
  proc497 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_63_o0 <= sig_64_o0;
      end if;
    end if;
  end process proc497;
  sig_64_o0 <= '1' when (sig_10_o0 = '1') else
               sig_65_o0;
  sig_65_o0 <= (sig_56_o0 or sig_66_o0);
  sig_66_o0 <= not(sig_67_o0);
  sig_67_o0 <= '0' when (sig_10_o0 = '1') else
               sig_61_o0;
  proc502 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_59_o0 <= sig_52_o0;
      end if;
    end if;
  end process proc502;
  sig_53_o0 <= (sig_13_o0 and sig_54_o0);
  proc504 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_54_o0 <= sig_55_o0;
      end if;
    end if;
  end process proc504;
  sig_55_o0 <= '1' when (sig_10_o0 = '1') else
               sig_56_o0;
  sig_56_o0 <= (sig_47_o0 or sig_57_o0);
  sig_57_o0 <= not(sig_58_o0);
  sig_58_o0 <= '0' when (sig_10_o0 = '1') else
               sig_52_o0;
  proc509 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_50_o0 <= sig_43_o0;
      end if;
    end if;
  end process proc509;
  sig_44_o0 <= (sig_13_o0 and sig_45_o0);
  proc511 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_45_o0 <= sig_46_o0;
      end if;
    end if;
  end process proc511;
  sig_46_o0 <= '1' when (sig_10_o0 = '1') else
               sig_47_o0;
  sig_47_o0 <= (sig_38_o0 or sig_48_o0);
  sig_48_o0 <= not(sig_49_o0);
  sig_49_o0 <= '0' when (sig_10_o0 = '1') else
               sig_43_o0;
  proc516 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_41_o0 <= sig_34_o0;
      end if;
    end if;
  end process proc516;
  sig_35_o0 <= (sig_13_o0 and sig_36_o0);
  proc518 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_36_o0 <= sig_37_o0;
      end if;
    end if;
  end process proc518;
  sig_37_o0 <= '1' when (sig_10_o0 = '1') else
               sig_38_o0;
  sig_38_o0 <= (sig_16_o0 or sig_39_o0);
  sig_39_o0 <= not(sig_40_o0);
  sig_40_o0 <= '0' when (sig_10_o0 = '1') else
               sig_34_o0;
  proc523 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_32_o0 <= sig_11_o0;
      end if;
    end if;
  end process proc523;
  sig_12_o0 <= (sig_13_o0 and sig_14_o0);
  proc525 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_14_o0 <= sig_15_o0;
      end if;
    end if;
  end process proc525;
  sig_15_o0 <= '1' when (sig_10_o0 = '1') else
               sig_16_o0;
  sig_16_o0 <= (sig_17_o0 or sig_31_o0);
  sig_31_o0 <= not(sig_9_o0);
  sig_17_o0 <= (sig_18_o0 or sig_23_o0);
  sig_23_o0 <= not(sig_24_o0);
  sig_24_o0 <= '0' when (sig_10_o0 = '1') else
               sig_25_o0;
  sig_25_o0 <= sig_30_o0 when (sig_26_o0 = '1') else
               sig_29_o0;
  proc533 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_30_o0 <= sig_11_o0;
      end if;
    end if;
  end process proc533;
  proc534 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_29_o0 <= sig_25_o0;
      end if;
    end if;
  end process proc534;
  sig_26_o0 <= (sig_13_o0 and sig_27_o0);
  proc536 : process(clk) is
  begin
    if rising_edge(clk) then
      if true then
        sig_27_o0 <= sig_28_o0;
      end if;
    end if;
  end process proc536;
  sig_28_o0 <= '1' when (sig_10_o0 = '1') else
               sig_17_o0;
  sig_18_o0 <= sig_19_o0(17);
  -- [("i0",16U,(20).o0),("i1",B,(21).o0),("i2",B,(22).o0)];
  sig_19_o0 <= sig_22_o0 & sig_21_o0 & sig_20_o0;
  sig_22_o0 <= out_ready;
  sig_21_o0 <= in_valid;
  sig_20_o0 <= in_x;
  sig_13_o0 <= not(sig_10_o0);
  sig_10_o0 <= reset;
  out_valid <= sig_2_o0;
  in_ready <= sig_269_o0;
  out_x <= sig_271_o0;
end architecture str;
